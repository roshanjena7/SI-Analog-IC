                                                                                                                                                                                               .PARAM vdd_var=1                                                                                                                                                                                                                                                                                                                                                                                                                      **Netlist                                                                                                                                                                                                          R1    vin     vout    1k                                                                                                                                                                                           C1    vout    GND     1p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 **Sources                                                                                                                                                                                                          vsin     vin     GND     0 PULSE(0 vdd_var 0.5n 1p 1p 20n)                                                                                                                                                                                                                                                                                                                                                                            **simulation                                                                                                                                                                                                       .OP                                                                                                                                                                                                                .TRAN 10p 40n                                                                                                                                                                                                                                                                                                                                                                                                                         .END                     
